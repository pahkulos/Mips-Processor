`define DELAY 20
module _32bit_alu_testbench(); 
reg   [31:0] inp_A,inp_B;
reg   [2:0] select;
wire  [31:0]out;

_32bit_alu alu32(out,inp_A,inp_B,select);
initial begin
//////////////////ADDER/////////////////////////
inp_A=32'b00000000000000000000000000000000; inp_B=32'b00000000000000000000000000000000; select=3'b000;
#`DELAY;
inp_A=32'b00000000000000000000000000000000; inp_B=32'b11111111111111111111111111111111; select=3'b000;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b00000000000000000000000000000000; select=3'b000;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b11111111111111111111111111111111; select=3'b000;
#`DELAY;

//////////////////XOR/////////////////////////
inp_A=32'b00000000000000000000000000000000; inp_B=32'b00000000000000000000000000000000; select=3'b001;
#`DELAY;
inp_A=32'b00000000000000000000000000000000; inp_B=32'b11111111111111111111111111111111; select=3'b001;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b00000000000000000000000000000000; select=3'b001;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b11111111111111111111111111111111; select=3'b001;
#`DELAY;


//////////////////SUB/////////////////////////
inp_A=32'b00000000000000000000000000000000; inp_B=32'b00000000000000000000000000000000; select=3'b010;
#`DELAY;
inp_A=32'b00000000000000000000000000000000; inp_B=32'b11111111111111111111111111111111; select=3'b010;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b00000000000000000000000000000000; select=3'b010;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b11111111111111111111111111111111; select=3'b010;
#`DELAY;

//////////////////SLT/////////////////////////
inp_A=32'b00000000000000000000000000000000; inp_B=32'b00000000000000000000000000000000; select=3'b100;
#`DELAY;
inp_A=32'b00000000000000000000000000000000; inp_B=32'b11111111111111111111111111111111; select=3'b100;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b00000000000000000000000000000000; select=3'b100;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b11111111111111111111111111111111; select=3'b100;
#`DELAY;

//////////////////NOR/////////////////////////
inp_A=32'b00000000000000000000000000000000; inp_B=32'b00000000000000000000000000000000; select=3'b101;
#`DELAY;
inp_A=32'b00000000000000000000000000000000; inp_B=32'b11111111111111111111111111111111; select=3'b101;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b00000000000000000000000000000000; select=3'b101;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b11111111111111111111111111111111; select=3'b101;
#`DELAY;

//////////////////AND/////////////////////////
inp_A=32'b00000000000000000000000000000000; inp_B=32'b00000000000000000000000000000000; select=3'b110;
#`DELAY;
inp_A=32'b00000000000000000000000000000000; inp_B=32'b11111111111111111111111111111111; select=3'b110;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b00000000000000000000000000000000; select=3'b110;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b11111111111111111111111111111111; select=3'b110;
#`DELAY;

//////////////////OR/////////////////////////
inp_A=32'b00000000000000000000000000000000; inp_B=32'b00000000000000000000000000000000; select=3'b111;
#`DELAY;
inp_A=32'b00000000000000000000000000000000; inp_B=32'b11111111111111111111111111111111; select=3'b111;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b00000000000000000000000000000000; select=3'b111;
#`DELAY;
inp_A=32'b11111111111111111111111111111111; inp_B=32'b11111111111111111111111111111111; select=3'b111;
#`DELAY;
end
 
 
initial
begin
$monitor("time = %2d, inp_A =%32b, inp_B=%32b, select=%3b, out=%32b", $time, inp_A, inp_B,select, out);
end
 
endmodule